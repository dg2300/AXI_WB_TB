//This is Testbench top
